// get data and sort 

// also outputs to the mux 
module ScoreBoardDisplay(); 
	


endmodule 