//sikender 


module ScoreBoard(); 


endmodule 