// ECE5440
// Sikender Shahid 1476
// Description: Access Control module compares 
// input passwords with stored password in the rom. 
// the comparator performs operation on 4bit values 
// with 4 entries in the ROM


