
`ifndef LCDController_vh
`define LCDController_vh

`define ENTER
`define USERID
`define PASSWORD
`define GAME
//A single HD44780U can display up to one 8-character line or two 8-character lines
