

module AccessControl_TEST_BENCH();

endmodule


